----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02.11.2023 23:38:55
-- Design Name: 
-- Module Name: libfram - package
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;


package libfram is
constant cnoCmd         : std_logic_vector(1 downto 0) := "00";
constant cFramReset     : std_logic_vector(1 downto 0) := "01";
constant cFramRead      : std_logic_vector(1 downto 0) := "10";
constant cFramWrite     : std_logic_vector(1 downto 0) := "11";
end libfram;

package body libfram is

end libfram;